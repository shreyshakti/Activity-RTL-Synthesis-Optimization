    Mac OS X            	   2       K                                      ATTR      K   �   �                  �   <  com.apple.quarantine    �   S  com.dropbox.attributes   q/0081;5cefecd6;Chrome;0E789C69-A87B-4A9B-AE8D-71038A4D5BB0 x��VJ)�/Hʯ�O��I�L���ON�Q�R�V�ML����%����RK��<�"���|W���L�b� ˀ@[[���Z Ȃe