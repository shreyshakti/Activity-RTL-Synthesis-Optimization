    Mac OS X            	   2  Q     �                                      ATTR      �   �   �                  �     com.apple.lastuseddate#PS       �   <  com.apple.quarantine   0   S  com.dropbox.attributes   ���\    k$9    q/0081;5cefecd6;Chrome;0E789C69-A87B-4A9B-AE8D-71038A4D5BB0 x��VJ)�/Hʯ�O��I�L���ON�Q�R�V�ML����%����RK���J��,�`�tgC�,s�R���r[[���Z �6�